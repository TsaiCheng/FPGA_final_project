module LED8x8(DATA_R,DATA_G,DATA_B,COMM,a,b,c,d,e,f,g,CLK,left,right,speed,rotation,clear,timeout);
	output reg[7:0] DATA_R,DATA_G,DATA_B;
	output reg[3:0] COMM;
	output reg a,b,c,d,e,f,g;
	input CLK,left,right,speed,rotation,clear,timeout;
	int test=0,origin=1,gg=0,score=0,rotationtime,find,fivetime=0,color=0,randomnum=0,n,n1,n2,n3;
	bit[7:0]one[7:0]=//正方型
		'{8'b11111111,
		8'b11111111,
		8'b11111111,
		8'b11111100,
		8'b11111100,
		8'b11111111,
		8'b11111111,
		8'b11111111};
	bit[7:0]two[7:0]=//一條線
		'{8'b11111111,
		8'b11111111,
		8'b11111110,
		8'b11111110,
		8'b11111110,
		8'b11111110,
		8'b11111111,
		8'b11111111};
	bit[7:0]three[7:0]=//左閃電
		'{8'b11111111,
		8'b11111111,
		8'b11111111,
		8'b11111101,
		8'b11111100,
		8'b11111110,
		8'b11111111,
		8'b11111111};
	bit[7:0]four[7:0]=//右閃電
		'{8'b11111111,
		8'b11111111,
		8'b11111110,
		8'b11111100,
		8'b11111101,
		8'b11111111,
		8'b11111111,
		8'b11111111};
	bit[7:0]five[7:0]=//左勺子
		'{8'b11111111,
		8'b11111111,
		8'b11111111,
		8'b11111110,
		8'b11111110,
		8'b11111100,
		8'b11111111,
		8'b11111111};
	bit[7:0]six[7:0]=//右勺子
		'{8'b11111111,
		8'b11111111,
		8'b11111100,
		8'b11111110,
		8'b11111110,
		8'b11111111,
		8'b11111111,
		8'b11111111};
	bit[7:0]seven[7:0]=//十字架
		'{8'b11111111,
		8'b11111111,
		8'b11111111,
		8'b11111110,
		8'b11111100,
		8'b11111110,
		8'b11111111,
		8'b11111111};
	bit[7:0]start[7:0]=//開始
		'{8'b01111110,
		8'b00000000,
		8'b01111110,
		8'b11111111,
		8'b00000000,
		8'b11110111,
		8'b11110111,
		8'b00000000};
	bit[7:0]zero[7:0]=//歸零
		'{8'b11111111,
		8'b11111111,
		8'b11111111,
		8'b11111111,
		8'b11111111,
		8'b11111111,
		8'b11111111,
		8'b11111111};
	bit[7:0]tmp[7:0];//暫存
	bit[7:0]now[7:0];//背景
	bit[7:0]R[7:0];
	bit[7:0]G[7:0];
	bit[7:0]B[7:0];
	bit[2:0] cnt,num;
	
	divfreq_1 (CLK_div_1,CLK);
	divfreq_2 (CLK_div_2,CLK);
	initial//初始化
		begin
		cnt=0;
		DATA_R=8'b11111111;
		DATA_G=8'b11111111;
		DATA_B=8'b11111111;
		COMM=4'b1000;
		end
	always @(posedge CLK_div_2)//下降
		begin
		if(clear==1)//歸零
			begin
			now=zero;
			R=zero;
			G=zero;
			B=zero;
			origin=1;
			gg=0;
			score=0;
			fivetime=0;
			end
		else
			for(n=0;n<=speed;++n)
				if(gg==0&&timeout==0)
					begin
					if(test==1||origin==1)//到底
						begin
						++fivetime;
						for(n1=0;n1<8;++n1)//檢查消掉
							begin
							test=0;
							for(n2=0;n2<8;++n2)
								if(now[n2][n1]==0)
									++test;
							if(test==8)//消掉
								begin
								++score;
								for(n2=7;n2>=0;--n2)
									for(n3=n1;n3>0;--n3)
										begin
										now[n2][n3]=now[n2][n3-1];
										R[n2][n3]=R[n2][n3-1];
										G[n2][n3]=G[n2][n3-1];
										B[n2][n3]=B[n2][n3-1];
										end
								for(n2=0;n2<8;++n2)
									begin
									now[n2][0]=1;
									R[n2][0]=1;
									G[n2][0]=1;
									B[n2][0]=1;
									end
								end
							end
						randomnum+=test;
						case(randomnum%7)//變換
							0:tmp=one;
							1:tmp=two;
							2:tmp=three;
							3:tmp=four;
							4:tmp=five;
							5:tmp=six;
							6:tmp=seven;
						endcase
						num=randomnum%7;
						++color;
						origin=0;
						rotationtime=0;
						end
					else//要繼續下降
						begin
						++fivetime;
						for(n1=0;n1<8;++n1)//now清掉tmp
							for(n2=0;n2<8;++n2)
								if(tmp[n1][n2]==0)
									begin
									now[n1][n2]=1;
									case(color%3)
										0:
											R[n1][n2]=1;
										1:
											G[n1][n2]=1;
										2:
											B[n1][n2]=1;
									endcase
									end
						if(fivetime%4==0)
							begin
							for(n1=7;n1>=0;--n1)//下降
								for(n2=7;n2>0;--n2)
									tmp[n1][n2]=tmp[n1][n2-1];
							for(n1=0;n1<8;++n1)//第一排歸零
								tmp[n1][0]=1;
							end
						end
					test=1;
					if(left==1)//左移
						begin
						randomnum+=2;
						for(n1=0;n1<8;++n1)
							if(tmp[0][n1]==0)
								begin
								test=0;
								break;
								end
						if(test==1)
							for(n1=1;n1<8;++n1)
								begin
								for(n2=0;n2<8;++n2)
									if(tmp[n1][n2]==0&&now[n1-1][n2]==0)
										begin
										test=0;
										break;
										end
								if(test==0)
									break;
								end
						if(test==1)
							begin
							for(n1=0;n1<7;++n1)
								for(n2=0;n2<8;++n2)
									tmp[n1][n2]=tmp[n1+1][n2];
							for(n1=0;n1<8;++n1)
								tmp[7][n1]=1;
							end
						end
					if(right==1)//右移
						begin
						randomnum+=1;
						for(n1=0;n1<8;++n1)
							if(tmp[7][n1]==0)
								begin
								test=0;
								break;
								end
						if(test==1)
							for(n1=0;n1<7;++n1)
								begin
								for(n2=0;n2<8;++n2)
									if(tmp[n1][n2]==0&&now[n1+1][n2]==0)
										begin
										test=0;
										break;
										end
								if(test==0)
									break;
								end
						if(test==1)
							begin
							for(n1=7;n1>0;--n1)
								for(n2=7;n2>=0;--n2)
									tmp[n1][n2]=tmp[n1-1][n2];
							for(n1=0;n1<8;++n1)
								tmp[0][n1]=1;
							end
						end
					/*if(rotation==1)//旋轉
							begin
							test=0;
							find=0;
							for(n1=0;n1<8;++n1)
								begin
								for(n2=0;n2<8;++n2)
									if(tmp[n1][n2]==0)
										begin
										find=1;
										case(num)
											1:
												case(rotationtime%2)
													0:
														if(n1<=4&&1<=n2&&n2<=5)
															if(now[n1+1][n2-1]==1&&now[n1+1][n2+1]==1&&now[n1+1][n2+2]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1+2][n2]=1;
																tmp[n1+3][n2]=1;
																tmp[n1+1][n2-1]=0;
																tmp[n1+1][n2+1]=0;
																tmp[n1+1][n2+2]=0;
																end
													1:
														if(1<=n1&&n1<=5&&n2<=4)
															if(now[n1-1][n2+1]==1&&now[n1+1][n2+1]==1&&now[n1+2][n2+1]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1][n2+2]=1;
																tmp[n1][n2+3]=1;
																tmp[n1-1][n2+1]=0;
																tmp[n1+1][n2+1]=0;
																tmp[n1+2][n2+1]=0;
																end
												endcase
											2:
												case(rotationtime%2)
													0:
														if(n1<=5&&1<=n2&&n2<=6)
															if(now[n1][n2+1]==1&&now[n1+1][n2-1]==1)
																begin
																test=1;
																tmp[n1+1][n2+1]=1;
																tmp[n1+2][n2+1]=1;
																tmp[n1][n2+1]=0;
																tmp[n1+1][n2-1]=0;
																end
													1:
														if(n1<=5&&1<=n2&&n2<=6)
															if(now[n1+1][n2+1]==1&&now[n1+2][n2+1]==1)
																begin
																test=1;
																tmp[n1][n2+1]=1;
																tmp[n1+1][n2-1]=1;
																tmp[n1+1][n2+1]=0;
																tmp[n1+2][n2+1]=0;
																end
												endcase
											3:
												case(rotationtime%2)
													0:
														if(n1<=5&&2<=n2)
															if(now[n1+1][n2-2]==1&&now[n1+2][n2]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1+1][n2]=1;
																tmp[n1+1][n2-2]=0;
																tmp[n1+2][n2]=0;
																end
													1:
														if(1<=n1&&n1<=6&&n2<=5)
															if(now[n1-1][n2+2]==1&&now[n1][n2+2]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1+1][n2+2]=1;
																tmp[n1-1][n2+2]=0;
																tmp[n1][n2+2]=0;
																end
												endcase
											4:
												case(rotationtime%4)
													0:
														if(n1<=5&&1<=n2&&n2<=6)
															if(now[n1][n2-1]==1&&now[n1+1][n2-1]==1&&now[n1+1][n2+1]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1][n2+1]=1;
																tmp[n1+2][n2]=1;
																tmp[n1][n2-1]=0;
																tmp[n1+1][n2-1]=0;
																tmp[n1+1][n2+1]=0;
																end
													1:
														if(n1<=5&&n2<=5)
															if(now[n1][n2+1]==1&&now[n1+2][n2]==1&&now[n1+2][n2+1]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1+1][n2]=1;
																tmp[n1+1][n2+2]=1;
																tmp[n1][n2+1]=0;
																tmp[n1+2][n2]=0;
																tmp[n1+2][n2+1]=0;
																end
													2:
														if(n1<=5&&1<=n2&&n2<=6)
															if(now[n1+1][n2-1]==1&&now[n1+1][n2+1]==1&&now[n1+2][n2+1]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1+2][n2-1]=1;
																tmp[n1+2][n2]=1;
																tmp[n1+1][n2-1]=0;
																tmp[n1+1][n2+1]=0;
																tmp[n1+2][n2+1]=0;
																end
													3:
														if(1<=n1&&n1<=6&&n2<=5)
															if(now[n1-1][n2+1]==1&&now[n1-1][n2+2]==1&&now[n1+1][n2+1]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1][n2+2]=1;
																tmp[n1+1][n2+2]=1;
																tmp[n1-1][n2+1]=0;
																tmp[n1-1][n2+2]=0;
																tmp[n1+1][n2+1]=0;
																end
												endcase
											5:
												case(rotationtime%4)
													0:
														if(n1<=5&&1<=n2&&n2<=6)
															if(now[n1+1][n2-1]==1&&now[n1+2][n2-1]==1&&now[n1+1][n2+1]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1+2][n2]=1;
																tmp[n1+2][n2+1]=1;
																tmp[n1+1][n2-1]=0;
																tmp[n1+2][n2-1]=0;
																tmp[n1+1][n2+1]=0;
																end
													1:
														if(1<=n1&&n1<=6&&n2<=5)
															if(now[n1-1][n2]==1&&now[n1-1][n2+1]==1&&now[n1+1][n2+1]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1+1][n2]=1;
																tmp[n1][n2+2]=1;
																tmp[n1-1][n2]=0;
																tmp[n1-1][n2+1]=0;
																tmp[n1+1][n2+1]=0;
																end
													2:
														if(n1<=5&&n2<=5)
															if(now[n1+1][n2]==1&&now[n1][n2+2]==1&&now[n1+1][n2+2]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1][n2+1]=1;
																tmp[n1+2][n2+1]=1;
																tmp[n1+1][n2]=0;
																tmp[n1][n2+2]=0;
																tmp[n1+1][n2+2]=0;
																end
													3:
														if(n1<=5&&2<=n2)
															if(now[n1][n2-1]==1&&now[n1+2][n2-1]==1&&now[n1+2][n2]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1+1][n2]=1;
																tmp[n1+1][n2-2]=1;
																tmp[n1][n2-1]=0;
																tmp[n1+2][n2-1]=0;
																tmp[n1+2][n2]=0;
																end
												endcase
											6:
												case(rotationtime%4)
													0:
														if(n1<=5&&1<=n2)
															if(now[n1+1][n2-1]==1)
																begin
																test=1;
																tmp[n1+2][n2]=1;
																tmp[n1+1][n2-1]=0;
																end
													1:
														if(n1<=5&&n2<=6)
															if(now[n1+2][n2]==1)
																begin
																test=1;
																tmp[n1+1][n2+1]=1;
																tmp[n1+2][n2]=0;
																end
													2:
														if(n1<=6&&n2<=6)
															if(now[n1+1][n2+1]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1+1][n2+1]=0;
																end
													3:
														if(1<=n1&&n2<=6)
															if(now[n1-1][n2+1]==1)
																begin
																test=1;
																tmp[n1][n2]=1;
																tmp[n1-1][n2+1]=0;
																end
												endcase
										endcase
										break;
										end
								if(test==1)
									++rotationtime;
								if(find==1)
									break;
								end
							end*/
					for(n1=0;n1<8;++n1)//檢查gg
						begin
						for(n2=0;n2<2;++n2)
							if(tmp[n1][n2]==0&&now[n1][n2]==0)
								begin
								gg=1;
								break;
								end
						if(gg==1)
							break;
						end
					if(gg==0)
						begin
						test=0;
						for(n1=7;n1>=0;--n1)//是否繼續下降
							begin
							for(n2=7;n2>=0;--n2)
								if(tmp[n2][n1]==0)
									begin
									if(n1==7)
										begin
										test=1;
										break;
										end
									else if(now[n2][n1+1]==0)
										begin
										test=1;
										break;
										end
									end
							if(test==1)
								break;
							end
						end
					for(n1=0;n1<8;++n1)//tmp丟到now
						for(n2=0;n2<8;++n2)
							if(tmp[n1][n2]==0)
								begin
								now[n1][n2]=0;
								case(color%3)
									0:
										R[n1][n2]=0;
									1:
										G[n1][n2]=0;
									2:
										B[n1][n2]=0;
								endcase
								end
					end
		end
	always @(posedge CLK_div_1)//顯示
		begin
		if(cnt>=7)
			cnt=0;
		else
			++cnt;
		COMM={1'b1,cnt};
		case(score)
			0:{a,b,c,d,e,f,g}=7'b0000001;
			1:{a,b,c,d,e,f,g}=7'b1001111;
			2:{a,b,c,d,e,f,g}=7'b0010010;
			3:{a,b,c,d,e,f,g}=7'b0000110;
			4:{a,b,c,d,e,f,g}=7'b1001100;
			5:{a,b,c,d,e,f,g}=7'b0100100;
			6:{a,b,c,d,e,f,g}=7'b0100000;
			7:{a,b,c,d,e,f,g}=7'b0001111;
			8:{a,b,c,d,e,f,g}=7'b0000000;
			9:{a,b,c,d,e,f,g}=7'b0000100;
		endcase
		if(origin==1||clear==1)//一開始
			begin
			DATA_R=start[cnt];
			DATA_G=8'b11111111;
			DATA_B=8'b11111111;
			end
		else
			begin
			DATA_R=R[cnt];
			DATA_G=G[cnt];
			DATA_B=B[cnt];
			end
		end
endmodule


module divfreq_1(output reg CLK_div,input CLK);
	reg[24:0] Count;
	
	always @(posedge CLK)
		begin
		if(Count>25000)
			begin
			Count<=25'b0;
			CLK_div<=~CLK_div;
			end
		else
			Count<=Count+1'b1;
		end
endmodule


module divfreq_2(output reg CLK_div,input CLK);
	reg[24:0] Count;
	
	always @(posedge CLK)
		begin
		if(Count>6250000)
			begin
			Count<=25'b0;
			CLK_div<=~CLK_div;
			end
		else
			Count<=Count+1'b1;
		end
endmodule
